// $Id: $
// File name:   input_sr.sv
// Created:     4/25/2016
// Author:      Dan Suciu
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: shift resgister for taking 8 bits and making d+ and d- for the input to the top level mapping
