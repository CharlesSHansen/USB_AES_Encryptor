mg101@ee215lnx07.ecn.purdue.edu.12627:1459956602