/home/ecegrid/a/mg101/ece337/USB_AES_Encryptor/source/USB_Reciever//pid_fifo.sv