/home/ecegrid/a/mg101/ece337/USB_AES_Encryptor/source/USB_Reciever//flex_stp_sr.sv