// $Id: $
// File name:   tb_usb_receiver.sv
// Created:     3/1/2016
// Author:      Charles Hansen
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: USB Receiver Testbench
