// $Id: $
// File name:   addRoundKey.sv
// Created:     4/24/2016
// Author:      Mitchel Bouma
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: add round key block

input addRoundKey();



endmodule